`timescale 1ns / 1ps
module tb_64x1_using_8x1_using_2x1();
reg [63:0]a;
reg [5:0]s;
wire y;
mux_64x1_using_8x1 g1(.y(y), .a(a), .s(s));
initial begin
s=6'b000000;a=64'b0;a[0]=1'b1;#5
s=6'b000001;a=64'b0;a[1]=1'b1;#5
s=6'b000010;a=64'b0;a[2]=1'b1;#5
s=6'b000011;a=64'b0;a[3]=1'b1;#5
s=6'b000100;a=64'b0;a[4]=1'b1;#5
s=6'b000101;a=64'b0;a[5]=1'b1;#5
s=6'b000110;a=64'b0;a[6]=1'b1;#5
s=6'b000111;a=64'b0;a[7]=1'b1;#5
s=6'b100100;a=64'b0;a[36]=1'b1;#5
s=6'b100110;a=64'b0;a[38]=1'b1;#5
s=6'b111100;a=64'b0;a[60]=1'b1;#5
s=6'b111101;a=64'b0;a[61]=1'b1;#5
s=6'b111110;a=64'b0;a[62]=1'b1;#5
s=6'b111111;a=64'b0;a[63]=1'b1;#5
$stop;
end
endmodule
