`timescale 1ns / 1ps
module tb_comparator();
reg [1:0]a,b;
wire [2:0]c;
comparator g1(.a(a), .b(b), .c(c));
initial begin
a[1]=0;a[0]=0;b[1]=0;b[0]=0;#5
a[1]=0;a[0]=0;b[1]=0;b[0]=1;#5
a[1]=0;a[0]=0;b[1]=1;b[0]=0;#5
a[1]=0;a[0]=0;b[1]=1;b[0]=1;#5
a[1]=0;a[0]=1;b[1]=0;b[0]=0;#5
a[1]=0;a[0]=1;b[1]=0;b[0]=1;#5
a[1]=0;a[0]=1;b[1]=1;b[0]=0;#5
a[1]=0;a[0]=1;b[1]=1;b[0]=1;#5
a[1]=1;a[0]=0;b[1]=0;b[0]=0;#5
a[1]=1;a[0]=0;b[1]=0;b[0]=1;#5
a[1]=1;a[0]=0;b[1]=1;b[0]=0;#5
a[1]=1;a[0]=0;b[1]=1;b[0]=1;#5
a[1]=1;a[0]=1;b[1]=0;b[0]=0;#5
a[1]=1;a[0]=1;b[1]=0;b[0]=1;#5
a[1]=1;a[0]=1;b[1]=1;b[0]=0;#5
a[1]=1;a[0]=1;b[1]=1;b[0]=1;#5
$stop;
end
endmodule
